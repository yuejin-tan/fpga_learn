-module ahb_epwm
-module ahb_lcd8080
-module ahb_null
-module ahb_seg7x8
-module ahb_sram
-module ahb_uart
-module AHBlite_Decoder
-module AHBlite_Interconnect
-module AHBlite_SlaveMUX
-module led_wf
-module top
-module PLL_FREQ
-topmoduleNum 2
-topmodule ahb_null
-topmodule top
