-module cm3_sys
-module top
-module PLL_25to200
-module led_wf
-module ahb_sram
-topmoduleNum 1
-topmodule top
