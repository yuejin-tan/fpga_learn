`timescale 1ns / 1ps 
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2024/03/16 10:31:59
// Design Name:
// Module Name: cm0_wrap
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module cm0_wrap(
    input wire clk,
    input wire RSTn,
    inout wire SWDIO,
    input wire SWCLK,

    //数码管接口
    output wire seg7_SH_CP,   //移位时钟
    output wire seg7_ST_CP,   //数据锁存时钟
    output wire seg7_DS,      //移位串行数据

    input wire RX_IN,
    output wire TX_OUT
  );

  //------------------------------------------------------------------------------
  // DEBUG IOBUF
  //------------------------------------------------------------------------------

  wire SWDO;
  wire SWDOEN;
  wire SWDI;

  assign SWDI = SWDIO;
  assign SWDIO = (SWDOEN) ? SWDO : 1'bz;

  // Interrupt

  wire [31: 0] IRQ;
  wire uartIntSig;
  /*Connect the IRQ with keyboard*/
  assign IRQ = {31'b0, uartIntSig};

  wire RXEV = 1'b0;

  // AHB

  wire [31: 0] HADDR;
  wire [ 2: 0] HBURST;
  wire HMASTLOCK;
  wire [ 3: 0] HPROT;
  wire [ 2: 0] HSIZE;
  wire [ 1: 0] HTRANS;
  wire [31: 0] HWDATA;
  wire HWRITE;
  wire [31: 0] HRDATA;
  wire HRESP;
  wire HMASTER;
  wire HREADY;

  // RESET AND DEBUG

  wire SYSRESETREQ;
  reg cpuresetn;

  always @(posedge clk or negedge RSTn)
    begin
      if (~RSTn)
        cpuresetn <= 1'b0;
      else if (SYSRESETREQ)
        cpuresetn <= 1'b0;
      else
        cpuresetn <= 1'b1;
    end

  wire CDBGPWRUPREQ;
  reg CDBGPWRUPACK;

  always @(posedge clk or negedge RSTn)
    begin
      if (~RSTn)
        CDBGPWRUPACK <= 1'b0;
      else
        CDBGPWRUPACK <= CDBGPWRUPREQ;
    end


  //------------------------------------------------------------------------------
  // Instantiate Cortex-M0 processor logic level
  //------------------------------------------------------------------------------
  parameter CODE_RAM_WIDTH = 14;
  parameter DATA_RAM_WIDTH = 12;

  cortexm0ds_logic u_logic (
                     // System inputs
                     .FCLK (clk),           //FREE running clock
                     .SCLK (clk),           //system clock
                     .HCLK (clk),           //AHB clock
                     .DCLK (clk),           //Debug clock
                     .PORESETn (RSTn),          //Power on reset
                     .HRESETn (cpuresetn),     //AHB and System reset
                     .DBGRESETn (RSTn),          //Debug Reset
                     .RSTBYPASS (1'b0),          //Reset bypass
                     .SE (1'b0),          // dummy scan enable port for synthesis

                     // Power management inputs
                     .SLEEPHOLDREQn (1'b1),          // Sleep extension request from PMU
                     .WICENREQ (1'b0),          // WIC enable request from PMU
                     .CDBGPWRUPACK (CDBGPWRUPACK),  // Debug Power Up ACK from PMU

                     // Power management outputs
                     .CDBGPWRUPREQ (CDBGPWRUPREQ),
                     .SYSRESETREQ (SYSRESETREQ),

                     // System bus
                     .HADDR (HADDR[31: 0]),
                     .HTRANS (HTRANS[1: 0]),
                     .HSIZE (HSIZE[2: 0]),
                     .HBURST (HBURST[2: 0]),
                     .HPROT (HPROT[3: 0]),
                     .HMASTER (HMASTER),
                     .HMASTLOCK (HMASTLOCK),
                     .HWRITE (HWRITE),
                     .HWDATA (HWDATA[31: 0]),
                     .HRDATA (HRDATA[31: 0]),
                     .HREADY (HREADY),
                     .HRESP (HRESP),

                     // Interrupts
                     .IRQ (IRQ),          //Interrupt
                     .NMI (1'b0),         //Watch dog interrupt
                     .IRQLATENCY (8'h0),
                     .ECOREVNUM (28'h0),

                     // Systick
                     .STCLKEN (1'b0),
                     .STCALIB (26'h0),

                     // Debug - JTAG or Serial wire
                     // Inputs
                     .nTRST (1'b1),
                     .SWDITMS (SWDI),
                     .SWCLKTCK (SWCLK),
                     .TDI (1'b0),
                     // Outputs
                     .SWDO (SWDO),
                     .SWDOEN (SWDOEN),

                     .DBGRESTART (1'b0),

                     // Event communication
                     .RXEV (RXEV),         // Generate event when a DMA operation completed.
                     .EDBGRQ (1'b0)          // multi-core synchronous halt request
                   );

  // AHBlite Interconncet
  wire HSEL_P0;
  wire [31: 0] HADDR_P0;
  wire [2: 0] HBURST_P0;
  wire HMASTLOCK_P0;
  wire [3: 0] HPROT_P0;
  wire [2: 0] HSIZE_P0;
  wire [1: 0] HTRANS_P0;
  wire [31: 0] HWDATA_P0;
  wire HWRITE_P0;
  wire HREADY_P0;
  wire HREADYOUT_P0;
  wire [31: 0] HRDATA_P0;
  wire HRESP_P0;

  wire HSEL_P1;
  wire [31: 0] HADDR_P1;
  wire [2: 0] HBURST_P1;
  wire HMASTLOCK_P1;
  wire [3: 0] HPROT_P1;
  wire [2: 0] HSIZE_P1;
  wire [1: 0] HTRANS_P1;
  wire [31: 0] HWDATA_P1;
  wire HWRITE_P1;
  wire HREADY_P1;
  wire HREADYOUT_P1;
  wire [31: 0] HRDATA_P1;
  wire HRESP_P1;

  wire HSEL_P2;
  wire [31: 0] HADDR_P2;
  wire [2: 0] HBURST_P2;
  wire HMASTLOCK_P2;
  wire [3: 0] HPROT_P2;
  wire [2: 0] HSIZE_P2;
  wire [1: 0] HTRANS_P2;
  wire [31: 0] HWDATA_P2;
  wire HWRITE_P2;
  wire HREADY_P2;
  wire HREADYOUT_P2;
  wire [31: 0] HRDATA_P2;
  wire HRESP_P2;

  wire HSEL_P3;
  wire [31: 0] HADDR_P3;
  wire [2: 0] HBURST_P3;
  wire HMASTLOCK_P3;
  wire [3: 0] HPROT_P3;
  wire [2: 0] HSIZE_P3;
  wire [1: 0] HTRANS_P3;
  wire [31: 0] HWDATA_P3;
  wire HWRITE_P3;
  wire HREADY_P3;
  wire HREADYOUT_P3;
  wire [31: 0] HRDATA_P3;
  wire HRESP_P3;

  AHBlite_Interconnect Interconncet(
                         .HCLK (clk),
                         .HRESETn (cpuresetn),

                         // CORE SIDE
                         .HADDR (HADDR),
                         .HTRANS (HTRANS),
                         .HSIZE (HSIZE),
                         .HBURST (HBURST),
                         .HPROT (HPROT),
                         .HMASTLOCK (HMASTLOCK),
                         .HWRITE (HWRITE),
                         .HWDATA (HWDATA),
                         .HRDATA (HRDATA),
                         .HREADY (HREADY),
                         .HRESP (HRESP),

                         // P0
                         .HSEL_P0 (HSEL_P0),
                         .HADDR_P0 (HADDR_P0),
                         .HBURST_P0 (HBURST_P0),
                         .HMASTLOCK_P0 (HMASTLOCK_P0),
                         .HPROT_P0 (HPROT_P0),
                         .HSIZE_P0 (HSIZE_P0),
                         .HTRANS_P0 (HTRANS_P0),
                         .HWDATA_P0 (HWDATA_P0),
                         .HWRITE_P0 (HWRITE_P0),
                         .HREADY_P0 (HREADY_P0),
                         .HREADYOUT_P0 (HREADYOUT_P0),
                         .HRDATA_P0 (HRDATA_P0),
                         .HRESP_P0 (HRESP_P0),

                         // P1
                         .HSEL_P1 (HSEL_P1),
                         .HADDR_P1 (HADDR_P1),
                         .HBURST_P1 (HBURST_P1),
                         .HMASTLOCK_P1 (HMASTLOCK_P1),
                         .HPROT_P1 (HPROT_P1),
                         .HSIZE_P1 (HSIZE_P1),
                         .HTRANS_P1 (HTRANS_P1),
                         .HWDATA_P1 (HWDATA_P1),
                         .HWRITE_P1 (HWRITE_P1),
                         .HREADY_P1 (HREADY_P1),
                         .HREADYOUT_P1 (HREADYOUT_P1),
                         .HRDATA_P1 (HRDATA_P1),
                         .HRESP_P1 (HRESP_P1),

                         // P2
                         .HSEL_P2 (HSEL_P2),
                         .HADDR_P2 (HADDR_P2),
                         .HBURST_P2 (HBURST_P2),
                         .HMASTLOCK_P2 (HMASTLOCK_P2),
                         .HPROT_P2 (HPROT_P2),
                         .HSIZE_P2 (HSIZE_P2),
                         .HTRANS_P2 (HTRANS_P2),
                         .HWDATA_P2 (HWDATA_P2),
                         .HWRITE_P2 (HWRITE_P2),
                         .HREADY_P2 (HREADY_P2),
                         .HREADYOUT_P2 (HREADYOUT_P2),
                         .HRDATA_P2 (HRDATA_P2),
                         .HRESP_P2 (HRESP_P2),

                         // P3
                         .HSEL_P3 (HSEL_P3),
                         .HADDR_P3 (HADDR_P3),
                         .HBURST_P3 (HBURST_P3),
                         .HMASTLOCK_P3 (HMASTLOCK_P3),
                         .HPROT_P3 (HPROT_P3),
                         .HSIZE_P3 (HSIZE_P3),
                         .HTRANS_P3 (HTRANS_P3),
                         .HWDATA_P3 (HWDATA_P3),
                         .HWRITE_P3 (HWRITE_P3),
                         .HREADY_P3 (HREADY_P3),
                         .HREADYOUT_P3 (HREADYOUT_P3),
                         .HRDATA_P3 (HRDATA_P3),
                         .HRESP_P3 (HRESP_P3)
                       );

  // AHB RAMCODE
  wire [CODE_RAM_WIDTH - 3: 0] RAMCODE_ADDR;
  wire [31: 0] RAMCODE_RDATA;
  wire [3: 0] RAMCODE_WREN;
  wire [31: 0] RAMCODE_WDATA;
  wire RAMCODE_CS;

  cmsdk_ahb_to_sram#(CODE_RAM_WIDTH) RAMCODE_Interface(
                     .HCLK (clk),
                     .HRESETn (cpuresetn),
                     .HSEL (HSEL_P0),
                     .HADDR (HADDR_P0[CODE_RAM_WIDTH - 1: 0]),
                     .HSIZE (HSIZE_P0),
                     .HTRANS (HTRANS_P0),
                     .HWDATA (HWDATA_P0),
                     .HWRITE (HWRITE_P0),
                     .HRDATA (HRDATA_P0),
                     .HREADY (HREADY_P0),
                     .HREADYOUT (HREADYOUT_P0),
                     .HRESP (HRESP_P0),

                     .SRAMRDATA (RAMCODE_RDATA),
                     .SRAMADDR (RAMCODE_ADDR),
                     .SRAMWEN (RAMCODE_WREN),
                     .SRAMWDATA (RAMCODE_WDATA),
                     .SRAMCS (RAMCODE_CS)
                   );

  cmsdk_fpga_sram#(CODE_RAM_WIDTH - 2) RAM_CODE(
                   .CLK (clk),
                   .RDATA (RAMCODE_RDATA),
                   .ADDR (RAMCODE_ADDR),
                   .WREN (RAMCODE_WREN),
                   .WDATA (RAMCODE_WDATA),
                   .CS (RAMCODE_CS)
                 );

  // AHB RAMDATA
  wire [DATA_RAM_WIDTH - 3: 0] RAMDATA_ADDR;
  wire [31: 0] RAMDATA_RDATA;
  wire [3: 0] RAMDATA_WREN;
  wire [31: 0] RAMDATA_WDATA;
  wire RAMDATA_CS;

  cmsdk_ahb_to_sram#(DATA_RAM_WIDTH) RAMDATA_Interface(
                     .HCLK (clk),
                     .HRESETn (cpuresetn),
                     .HSEL (HSEL_P1),
                     .HADDR (HADDR_P1[DATA_RAM_WIDTH - 1: 0]),
                     .HSIZE (HSIZE_P1),
                     .HTRANS (HTRANS_P1),
                     .HWDATA (HWDATA_P1),
                     .HWRITE (HWRITE_P1),
                     .HRDATA (HRDATA_P1),
                     .HREADY (HREADY_P1),
                     .HREADYOUT (HREADYOUT_P1),
                     .HRESP (HRESP_P1),

                     .SRAMRDATA (RAMDATA_RDATA),
                     .SRAMADDR (RAMDATA_ADDR),
                     .SRAMWEN (RAMDATA_WREN),
                     .SRAMWDATA (RAMDATA_WDATA),
                     .SRAMCS (RAMDATA_CS)
                   );

  cmsdk_fpga_sram#(DATA_RAM_WIDTH - 2) RAM_DATA(
                   .CLK (clk),
                   .RDATA (RAMDATA_RDATA),
                   .ADDR (RAMDATA_ADDR),
                   .WREN (RAMDATA_WREN),
                   .WDATA (RAMDATA_WDATA),
                   .CS (RAMDATA_CS)
                 );

  // uart
  ahb_uart ahb_uart1(
             .HCLK ( clk ),
             .HRESETn ( cpuresetn ),

             .HSEL ( HSEL_P2 ),
             .HADDR ( HADDR_P2[ 15: 0 ] ),
             .HTRANS ( HTRANS_P2 ),
             .HSIZE ( HSIZE_P2 ),
             .HWRITE ( HWRITE_P2 ),
             .HWDATA ( HRDATA_P2 ),
             .HREADY ( HREADY_P2 ),

             .HREADYOUT ( HREADYOUT_P2 ),
             .HRDATA ( HRDATA_P2 ),
             .HRESP ( HRESP_P2 ),

             .INT_REQ( uartIntSig ),
             .TX_OUT( TX_OUT ),
             .RX_IN( RX_IN)
           );

  //  SEG7
  ahb_seg7x8 seg_inst(
               .HCLK ( clk ), //时钟
               .HRESETn ( cpuresetn ), //复位

               .HSEL ( HSEL_P3 ), // AHB inputs，设备选择
               .HADDR ( HADDR_P3[ 15: 0 ] ), //地址
               .HTRANS ( HTRANS_P3 ), //传输控制信号
               .HSIZE ( HSIZE_P3 ),  //传输大小
               .HWRITE ( HWRITE_P3 ), //写控制
               .HWDATA ( HRDATA_P3 ), //写数据
               .HREADY ( HREADY_P3 ), //传输完成

               .HREADYOUT ( HREADYOUT_P3 ), // AHB Outputs，设备准备信号
               .HRDATA ( HRDATA_P3 ), //读取到的数据
               .HRESP ( HRESP_P3 ), //设备响应

               .SH_CLK( seg7_SH_CP ),
               .LD_CLK( seg7_ST_CP ),
               .HC_DAT( seg7_DS)
             );

endmodule
